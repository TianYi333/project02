----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 2023/09/01 09:19:03
-- Design Name: 
-- Module Name: fun_servo - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package bus_multiplexer_pkg is
    type bus_array is array(natural range <>) of std_logic_vector(31 downto 0);
end package;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use work.bus_multiplexer_pkg.all;

Library xpm;
use xpm.vcomponents.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity fun_servo is
    generic(
        async_en        : std_logic:='0';
        regs_num        : integer:=17;
        runtime_num     : std_logic_vector(31 downto 0):=X"0773_5940"  -- 1s in 125MHz
    );
    Port (
        gtx_clk     		        : in  std_logic;
        rst                         : in  std_logic;
        -- rx cmd data
        rx_data_valid               : in  std_logic;
        rx_data_last                : in  std_logic;
        rx_data_data                : in  std_logic_vector(7 downto 0);
        -- tx data
        tx_data_valid               : out std_logic:='0';
        tx_data_last                : out std_logic:='0';
        tx_data_data                : out std_logic_vector(7 downto 0):=(others => '0');
        ini_status                  : out std_logic_Vector(3 downto 0):=(others => '0');
        -- angle servo
        angle_servo                 : out std_logic_Vector(15 downto 0):=(others => '0');
        -- uart
        UART_DIR                    : out   std_logic:='0';
        UART_IO                     : inout    std_logic
    );
end fun_servo;

architecture Behavioral of fun_servo is
    signal    ini_status1                :  std_logic_vector(3 downto 0):=(others => '0');
    
    signal    tx_data_last1              :  std_logic:='0';
    signal    angle_servo1                 : std_logic_Vector(15 downto 0):=(others => '0');
    -- uart io
    signal  uart_rx     : std_logic:='0';
    signal  uart_rx1     : std_logic:='0';
    signal  uart_tx     : std_logic:='0';
    signal  uart_ctrl   : std_logic:='Z';

    component UART
        Port (
            clk_in                : in    std_logic;
            UART_RX               : in    std_logic;
            UART_TX               : out   std_logic:='1';
            UART_DATA_IN_READY    : out   std_logic:='0';
            UART_DATA_IN          : in    std_logic_vector (7 downto 0);
            UART_DATA_IN_VALID    : IN    std_logic ;
            UART_DATA_OUT_END     : OUT   std_logic:='0';
            UART_DATA_OUT         : OUT   std_logic_vector (7 downto 0);
            UART_DATA_OUT_VALID   : OUT   STD_LOGIC
        );
    end component;

    signal  UART_DATA_IN_READY     :     std_logic:='0';
    signal  UART_DATA_OUT          :     std_logic_vector (7 downto 0);
    signal  UART_DATA_OUT_VALID    :     std_logic ;
    signal  UART_DATA_OUT_END      :     std_logic;

    component servo_tx
        generic(
            tx_head_01             : std_logic_vector(7 downto 0):=X"12";
            tx_head_02             : std_logic_vector(7 downto 0):=X"4C"
        );
        Port (
            aclk                      : in std_logic;
            rst                       : in std_logic;
            tx_data_in                : in std_logic_vector(7 downto 0);
            tx_data_in_valid          : in std_logic;
            servo_id                  : in std_logic_vector(7 downto 0);
            UART_DATA_IN_READY        : in std_logic;
            tx_data_out               : out std_logic_vector(7 downto 0);
            tx_data_out_valid         : out std_logic;
            tx_data_out_end           : out std_logic:='0'
        );
    end component;

    signal        tx_data_in                :  std_logic_vector(7 downto 0);
    signal        tx_data_in_valid          :  std_logic;
    signal        tx_servo_id               :  std_logic_vector(7 downto 0):=(others => '0');
    signal        tx_data_out               :  std_logic_vector(7 downto 0);
    signal        tx_data_out_valid         :  std_logic:='0';
    signal        tx_data_out_end           :  std_logic:='0';
    signal        tx_data_out_end1          :  std_logic:='0';

    component servo_rx
        Port (
            aclk                      : in std_logic;
            rst                       : in std_logic;
            rx_data_in                : in std_logic_vector(7 downto 0);
            rx_data_in_valid          : in std_logic;
            servo_id                  : in std_logic_vector(7 downto 0);
            error_code                : out std_logic_vector(7 downto 0):=(others => '0');
            rx_data_out               : out std_logic_vector(7 downto 0):=(others => '0');
            rx_data_out_valid         : out std_logic:='0';
            rx_data_out_last          : out std_logic:='0'
        );
    end component;

    signal        rx_data_in                :  std_logic_vector(7 downto 0);
    signal        rx_data_in_valid          :  std_logic;
    signal        error_code                :  std_logic_vector(7 downto 0):=(others => '0');
    signal        rx_servo_id               :  std_logic_vector(7 downto 0):=(others => '0');
    signal        rx_data_out               :  std_logic_vector(7 downto 0):=(others => '0');
    signal        rx_data_out_valid         :  std_logic:='0';
    signal        rx_data_out_last          :  std_logic:='0';

    signal        state_fun_servo           : std_logic_vector(3 downto 0):=(others => '1');        -- ��ʼ��״̬��ΪF
    signal        state_send_reg            : std_logic_vector(3 downto 0):=(others => '0');
    signal        length_reg                : std_logic_vector(3 downto 0):=(others => '0');
    signal        length_cnt                : std_logic_vector(3 downto 0):=(others => '0');

    signal  rx_data_valid1  : std_logic:='0';
    signal  runtime_cnt     : std_logic_Vector(31 downto 0):=(others => '0');

    signal  state_output_angle      : std_logic_vector(3 downto 0):=(others => '0');
    
    type ini_array  is array(0 to 10) of std_logic_vector(7 downto 0);
    signal  read_angle      : ini_array:=(
    0 => X"0A",     -- ���Ƕ�
    1 => X"02",     -- ���ݳ���
                    -- ����ʵ��Ϊ0
    others => (others => '0')
    );
    
    signal  read_angle_index       : integer:=0;       -- ���Ƕ�ʱ���ڷ������ݼ���
    signal  read_error_cnt          : integer:=0;       -- ���Ƕ�ʧ�ܣ�
    signal  send_angle      : ini_array:=(
    0 => X"08",     -- д�Ƕ�
    1 => X"07",     -- ���ݳ���
    2 => X"00",     -- ID
    3 => X"00",     -- �Ƕȵ�8λ    -- ʵ��ʹ��angle_servo1����
    4 => X"00",     -- �Ƕȸ�8λ 
    5 => X"E8",     -- ʱ���8λ 
    6 => X"03",     -- ʱ���8λ    -- ʱ�䶨Ϊ1s
    7 => X"00",     -- ���ʵ�8λ 
    8 => X"00",     -- ���ʸ�8λ 
    others => (others => '0')
    );
    signal  send_angle_index       : integer:=0;       -- д�Ƕ�ʱ���ڷ������ݼ���

--COMPONENT ila_0

--PORT (
--	clk : IN STD_LOGIC;



--	probe0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0); 
--	probe1 : IN STD_LOGIC_VECTOR(7 DOWNTO 0); 
--	probe2 : IN STD_LOGIC_VECTOR(0 DOWNTO 0); 
--	probe3 : IN STD_LOGIC_VECTOR(0 DOWNTO 0); 
--	probe4 : IN STD_LOGIC_VECTOR(7 DOWNTO 0); 
--	probe5 : IN STD_LOGIC_VECTOR(0 DOWNTO 0); 
--	probe6 : IN STD_LOGIC_VECTOR(7 DOWNTO 0); 
--	probe7 : IN STD_LOGIC_VECTOR(0 DOWNTO 0); 
--	probe8 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
--	probe9 : IN STD_LOGIC_VECTOR(0 DOWNTO 0)
--);
--END COMPONENT  ;

    
begin

--isnt_ila0 : ila_0
--PORT MAP (
--	clk => gtx_clk,



--	probe0 => state_fun_servo, 
--	probe1 => rx_data_out, 
--	probe2(0) => rx_data_out_valid,
--	probe3(0) => rx_data_out_last,
--	probe4 => rx_data_in,
--	probe5(0) => rx_data_in_valid,
--	probe6 => tx_data_out,
--	probe7(0) => tx_data_out_valid,
--	probe8(0) => UART_RX,
--	probe9(0) => uart_ctrl
	
--);

    tx_data_last <= tx_data_last1;
    main_state_gen : process(gtx_clk)
    begin
        if rising_edge(gtx_clk) then
--            ini_status1 <= '0';
            rx_data_valid1 <= rx_data_valid;
            tx_data_out_end1 <= tx_data_out_end;
--            if rst = '1'    then
--                state_fun_servo <= (others => '0');
--            else
                case    state_fun_servo is
                    when    X"0"    =>      -- �յ���λ����Ϣ�����͸�servo                        
                        if rx_data_valid = '1'  then
                            length_reg <= length_reg + '1';
                            tx_data_in <= rx_data_data;
                            tx_data_in_valid <= '1';
                            uart_ctrl <= '0';
                            if rx_data_valid1 = '0' then
                                tx_servo_id <= rx_data_data;
                                rx_servo_id <= rx_data_data;
                            end if;
                            if rx_data_last = '1'  then
                                state_fun_servo <= state_fun_servo + '1';
                            end if;
                        else
                            length_reg <= (others => '0');
                            tx_data_in_valid <= '0';
                            uart_ctrl <= 'Z';
                        end if;
                    when    X"1"    =>
                        state_fun_servo <= state_fun_servo + '1';
                        tx_data_in <= (others => '0');
                        tx_data_in_valid <= '0';
                    when    X"2"    =>  -- �ȴ�tx_data_out_end
                        if tx_data_out_end1 = '0' and tx_data_out_end = '1' then
                            state_fun_servo <= state_fun_servo + '1';
                        end if;
                    when    X"3"    =>  -- �ȴ� UART_DATA_IN_READY
                        if UART_DATA_IN_READY = '1' then
                            state_fun_servo <= state_fun_servo + '1';
                            runtime_cnt <= (others => '0');
                        end if;
                    when    X"4"    =>  -- ׼������servo���ݲ����͸���λ��
                        uart_ctrl <= '1';
                        tx_data_data  <= rx_data_out;
                        tx_data_valid <= rx_data_out_valid;
                        tx_data_last1  <=  rx_data_out_last;
                        if tx_data_last1 = '1' and rx_data_out_last = '0' then
                            state_fun_servo <= state_fun_servo + '1';
                        else
                            runtime_cnt <= runtime_cnt + '1';
                            if runtime_cnt = runtime_num    then
                                state_fun_servo <= X"6";
                            end if;
                        end if;
                    when    X"5"    =>
                        tx_data_last1 <= '0';
                        tx_data_data <= (others => '0');
                        tx_data_valid <= '0';
                        state_fun_servo <= (others => '0');
                    when    X"6"    =>
                        tx_data_data <= (others => '1');
                        tx_data_valid <= '1';
                        state_fun_servo <= state_fun_servo + '1';
                    when    X"7"    =>      -- rx time error
                        tx_data_data <= (others => '1');
                        tx_data_valid <= '1';
                        state_fun_servo <= state_fun_servo + '1';
                    when    X"8"    =>
                        tx_data_data <= (others => '1');
                        tx_data_valid <= '1';
                        state_fun_servo <= state_fun_servo + '1';
                    when    X"9"    =>
                        tx_data_data <= (others => '1');
                        tx_data_valid <= '1';
                        tx_data_last1 <= '1';
                        state_fun_servo <= state_fun_servo + '1';
                    when    X"A"    =>
                        tx_data_data <= (others => '0');
                        tx_data_valid <= '0';
                        tx_data_last1 <= '0';
                        state_fun_servo <= (others => '0');
                    -----------------------------------------------------------------
                    -- ini state+   20240224
                    when    X"B"    =>
                        tx_data_in_valid <= '0';
                        if tx_data_out_end1 = '0' and tx_data_out_end = '1' then
                            state_fun_servo <= X"E";
                        end if;
                    when    X"C"    =>   -- ��ɳ�ʼ��
                        if UART_DATA_IN_READY = '1' then
                            state_fun_servo <= X"0"; 
                            uart_ctrl <= '1';    
                            ini_status <= X"1";                       
                        end if;                        
                    when    X"D"    =>   -- ���ͽǶ�
                        if send_angle_index = 10 then
                            state_fun_servo <= X"C";
                            tx_data_in_valid <= '0';
                        else
                            uart_ctrl <= '0';
                            tx_data_in_valid <= '1';
                            send_angle_index <= send_angle_index + 1;                            
                            case send_angle_index is
                                when    3   =>
                                    tx_data_in <= angle_servo1(7 downto 0);
                                when    4   =>
                                    tx_data_in <= angle_servo1(15 downto 8);
                                when    others  =>
                                    tx_data_in <= send_angle(send_angle_index);
                            end case;
                        end if;
                    when    X"E"    =>   -- ׼�����սǶ�                           
                        if UART_DATA_IN_READY = '1' then
                            uart_ctrl <= '1';                            
                        end if;
                        if rx_data_out_last = '1' then
                            state_fun_servo <= X"D";
                        else
                            runtime_cnt <= runtime_cnt + '1';
                            if runtime_cnt = runtime_num    then
--                            if runtime_cnt = X"0000_f010"    then     --sim
                                state_fun_servo <= X"F";
                            end if;
                        end if;                      
                    when    X"F"    =>      -- ���Ƕ�
                        rx_servo_id <= read_angle(0);
                        runtime_cnt <= (others => '0');
                        if read_error_cnt = 10 then
                            ini_status <= X"F";
                            state_fun_servo <= X"0";
                        else
                            uart_ctrl <= '0';
                            tx_data_in_valid <= '1';
                            tx_data_in <= read_angle(read_angle_index);
                            if read_angle_index < 10 then
                                read_angle_index <= read_angle_index + 1;
                            else
                                read_angle_index <= 0;
                                state_fun_servo <= X"B";
                                read_error_cnt <= read_error_cnt + 1;
                            end if;
                        end if;
                    when    others  =>
                        state_fun_servo <= (others => '0');
                end case;
            end if;
--        end if;
    end process;

    inst_uart_io : IOBUF
        generic map (
            DRIVE => 12,
            IOSTANDARD => "DEFAULT",
            SLEW => "SLOW")
        port map (
            O => uart_rx1,     -- Buffer output
            IO => UART_IO,   -- Buffer inout port (connect directly to top-level port)
            I => uart_tx,     -- Buffer input
            T => uart_ctrl      -- 3-state enable input, high=input, low=output 
        );
    uart_rx <= uart_rx1 when uart_ctrl = '1' else '1';
    UART_DIR <= uart_ctrl;


    inst_servo_UART : UART
        port map(
            clk_in                  =>  gtx_clk             ,
            UART_RX                 =>  UART_RX            ,
            UART_TX                 =>  UART_TX            ,
            UART_DATA_IN_READY      =>  UART_DATA_IN_READY ,
            UART_DATA_IN            =>  tx_data_out       ,
            UART_DATA_IN_VALID      =>  tx_data_out_valid ,
            UART_DATA_OUT_END       =>  UART_DATA_OUT_END  ,
            UART_DATA_OUT           =>  UART_DATA_OUT      ,
            UART_DATA_OUT_VALID     =>  UART_DATA_OUT_VALID
        );

    inst_servo_tx : servo_tx
        port map(
            aclk                    =>  gtx_clk           ,
            rst                     =>  rst               ,
            tx_data_in              =>  tx_data_in        ,
            tx_data_in_valid        =>  tx_data_in_valid  ,
            servo_id                =>  tx_servo_id       ,
            UART_DATA_IN_READY      =>  UART_DATA_IN_READY,
            tx_data_out             =>  tx_data_out       ,
            tx_data_out_valid       =>  tx_data_out_valid,
            tx_data_out_end         =>  tx_data_out_end
        );

    rx_data_in <= UART_DATA_OUT;
    rx_data_in_valid <= UART_DATA_OUT_VALID;

    inst_servo_rx : servo_rx
        port map(
            aclk                    =>  gtx_clk          ,
            rst                     =>  rst              ,
            rx_data_in              =>  rx_data_in       ,
            rx_data_in_valid        =>  rx_data_in_valid ,
            servo_id                =>  rx_servo_id      ,
            error_code              =>  error_code       ,
            rx_data_out             =>  rx_data_out      ,
            rx_data_out_valid       =>  rx_data_out_valid,
            rx_data_out_last        =>  rx_data_out_last
        );

    process(gtx_clk)
    begin
        if rising_edge(gtx_clk) then
            case    state_output_angle  is
                when    X"0"    =>
                    if tx_data_out_valid = '1' and  tx_data_out = X"12" then
                        state_output_angle <= state_output_angle + '1';
                    end if;
                when    X"1"    =>
                    if tx_data_out_valid = '1'   then
                        if tx_data_out = X"4C" then
                            state_output_angle <= state_output_angle + '1';
                        else
                            state_output_angle <= X"0";
                        end if;
                    end if;
                when    X"2"    =>
                    if tx_data_out_valid = '1'   then
                        if tx_data_out = X"0A" then
                            state_output_angle <= state_output_angle + '1';
                        else
                            state_output_angle <= X"0";
                        end if;
                    end if;
                when    X"3"    =>
                    if tx_data_out_valid = '1'   then
--                        if tx_data_out = X"01" then
                            state_output_angle <= state_output_angle + '1';
--                        else
--                            state_output_angle <= X"0";
--                        end if;
                    end if;
                when    X"4"    =>
                    if rx_data_out_valid = '1'  then
                        if rx_data_out = X"0A" then
                            state_output_angle <= state_output_angle + '1';
                        else
                            state_output_angle <= X"0";
                        end if;
                    end if;
                when    X"5"    =>
                    if rx_data_out_valid = '1'  then
                        if rx_data_out = X"03" then
                            state_output_angle <= state_output_angle + '1';
                        else
                            state_output_angle <= X"0";
                        end if;
                    end if;
                when    X"6"    =>
                    if rx_data_out_valid = '1' then
                        state_output_angle <= state_output_angle + '1';
                    end if;
                when    X"7"    =>
                    if rx_data_out_valid = '1' then
                        angle_servo1(7 downto 0) <= rx_data_out;
                        state_output_angle <= state_output_angle + '1';
                    end if;
                when    X"8"    =>
                    if rx_data_out_valid = '1' then
                        angle_servo1(15 downto 8) <= rx_data_out;
                        state_output_angle <= X"0";
                    end if;
                when    others  =>

            end case;
        end if;
    end process;
angle_servo <= angle_servo1;
end Behavioral;
